LIBRARY ieee;
USE ieee.std_logic_1164.all;

PACKAGE display7seg_package IS
	COMPONENT display7seg IS
		PORT(num : IN std_logic_vector(3 DOWNTO 0);
			seg1 : OUT std_logic_vector(6 DOWNTO 0));
	END COMPONENT;
END display7seg_package;